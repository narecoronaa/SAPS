* AC Analysis, 1.2k lowPass, 2nd order Chebyshev 0.08 dB, 1 stage using AD8657

* Input signal for AC and transient sinusoidal analysis
VIN IN 0 AC 1 DC 0 SINE(0 4.94 118)
* VNOISE IN 0 AC 0 DC 0

XA IN OUT VCCG VEEG 0 multipleFeedbacklowPassStageA

VP VCCG 0 5
VM VEEG 0 -5

*Simulation directive lines for AC Analysis
.AC DEC 100 120 40k
*.TRAN 1n 3.29m
*.NOISE V(OUT) VNOISE DEC 100 120 40k
.SUBCKT multipleFeedbacklowPassStageA IN OUT VCC VEE GND
X1 GND INM VCC VEE OUT AD8657
R1 IN 1 100k
R2 1 INM 47k
R5 1 OUT 100k
C1 1 GND 4.7n
C2 INM OUT 1n
.ENDS multipleFeedbacklowPassStageA

* AD8657 SPICE Macro-model Typical Values
* Description: Amplifier
* Generic Desc: 3/18V, CMOS, OP, Low Pwr, RRIO, 2X
* Developed by: VW ADSJ
* Revision History: 08/10/2012 - Updated to new header style
* 1.1 (01/2011)
* Copyright 2010, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: VSY=18V, T=25�C
*
* END Notes
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT AD8657          1   2   99  50  45
*
* INPUT STAGE
*
M1   4  7  8  8 PIX L= 1.000E-06 W= 1.532E-04
M2   6  2  8  8 PIX L= 1.000E-06 W=1.532E-04
M3  14  7 18 18 NIX L=1.000E-06 W=4.085E-04
M4  16  2 18 18 NIX L=1.000E-06 W=4.085E-04
RD1  4 50 2.0E+04
RD2  6 50 2.0E+04
RD3 99 14 2.0E+04
RD4 99 16 2.0E+04
C1   4  6 9.4750E-12
C2  14 16 9.4750E-12
I1  99  8 1.722E-05
I2  18 50 1.722E-05
V1  99  9 1.429E-01
V2  19 50 1.429E-01
D1   8  9 DX
D2  19 18 DX
EOS  7  1 POLY(4) (73,98) (22,98) (81,98) (83,98) 3.500E-04 1 1 1 1
IOS  1  2 2.000E-11
CDiff  1 2 3.5E-12
Cin1   1 50 10.5E-12
Cin2   2 50 10.5E-12
*
*
* CMRR
*
E1  72 98 POLY(2) (1,98) (2,98) 0 6.817E-02 6.817E-02
R10 72 73 2.894E+02
R20 73 98 1.592E-02
C10 72 73 1.000E-06
*
* PSRR
*
EPSY 21 98 POLY(1) (99,50) -1.757E+02 9.762E+00
RPS1 21 22 3.183E+03
RPS2 22 98 7.958E-01
CPS1 21 22 1.000E-06
*
* VOLTAGE NOISE 
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 4.5165E+01
RN2 81 98 1
*
* FLICKER NOISE 
*
DFN 82 98 DNOISE
VFN 82 98 DC 0.6551
HFN 83 98 POLY(1) VFN 1.000E-03 1.000E+00
RFN 83 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) -1.74975E-05 5.031E-08
EVP  97 98 POLY(1) (99,50) -1.05 0.25
EVN  51 98 POLY(1) (50,99) 1.45 0.3

*
* GAIN STAGE
*
G1 98 30 POLY(2) (4,6) (14,16) 0 5.693E-05 5.693E-05
R1 30 98 1.000E+06
RZ 30 31 8.2720E+03
CF 45 31 5.60E-10
D3 30 97 DX
D4 51 30 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L= 2.000E-06 W=2.450E-04
M6  45 47 50 50 NOX L= 2.000E-06 W=1.591E-04
EG1 99 46 POLY(1) (98,30) 3.347E-01 1
EG2 47 50 POLY(1) (30,98) 3.216E-01 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=1.000E-05,VTO=-0.3,LAMBDA=0.01,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=4.000E-05,VTO=+0.3,LAMBDA=0.01,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=4.000E-05,VTO=-0.5,LAMBDA=0.01)
.MODEL NIX NMOS (LEVEL=2,KP=1.500E-05,VTO=0.5,LAMBDA=0.01)
.MODEL DX D(IS=1E-14,RS=0.1)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=1.5E-10)
*
*
.ENDS AD8657
*
*$





